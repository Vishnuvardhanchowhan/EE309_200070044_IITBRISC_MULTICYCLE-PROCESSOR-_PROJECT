library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
use ieee.math_real.all;

library work;
use work.basic.all;

entity IITB_RISC is
	port(clk,reset: in std_logic;
			clock_50: in bit;
			r0      : out std_logic_vector(15 downto 0);
		   r1      : out std_logic_vector(15 downto 0);
   		r2      : out std_logic_vector(15 downto 0);
	   	r3      : out std_logic_vector(15 downto 0);
		   r4      : out std_logic_vector(15 downto 0);
		   r5      : out std_logic_vector(15 downto 0);
		   r6      : out std_logic_vector(15 downto 0);
		   r7      : out std_logic_vector(15 downto 0));
end entity;

architecture behave of IITB_RISC is
	signal	m_mem_a       :   std_logic;
	signal	m_a3_0,m_a3_1 :   std_logic;
	signal	m_d3_0,m_d3_1 :   std_logic;
	signal	m_z           :   std_logic;
	signal m_comp_a,m_comp_b : std_logic;
	signal	m_op2_0,m_op2_1	        :   std_logic;
	signal	wr_mem        :   std_logic;   --write on memory
	signal	rd_mem        :   std_logic;   --read memory
	signal	wr_rf         :   std_logic;   --write on register file
	signal   m_a2			  :  std_logic;
	signal   m_op1_0,m_op1_1         :  std_logic;
	-----enable---------------------
	signal	en_ir,en_irf        :   std_logic;  --enable instruction register
	signal   en_A   : std_logic;
	signal	en_c,en_z     :   std_logic;
	signal	op_sel        :   std_logic;   --operation select by alu
	signal	condition_code:  std_logic_vector(1 downto 0);    --last 2 bits of IR
	signal	equ      :  std_logic;  --comparator
	signal	C,Z      :  std_logic;  --carry,zero
	signal	op_code  :  std_logic_vector(3 downto 0);  --first 4 bits of IR which is op_code
begin
	datapath_risc : datapath
			port map(
		m_mem_a	       => m_mem_a,
		m_a3_0         => m_a3_0,
		m_a3_1 	       => m_a3_1,
		m_d3_0         => m_d3_0,
		m_d3_1 	       => m_d3_1,
		m_z            => m_z,
		m_op2_0	       => m_op2_0,
		m_op2_1	       => m_op2_1,
		m_a2          => m_a2,
		m_op1_0          => m_op1_0,
		m_op1_1          => m_op1_1,
		wr_mem         => wr_mem,  
		rd_mem         => rd_mem,  
		wr_rf          => wr_rf,   
		en_ir          => en_ir,   
		en_irf      => en_irf, 
		en_A           => en_A,  
		en_c           => en_c,
		m_comp_a       => m_comp_a,
		m_comp_b       => m_comp_b,
		en_z           => en_z,
		op_sel         => op_sel,   
		equ            => equ,    
		C              => C,
		Z              => Z,  
		op_code        => op_code,
		condition_code => condition_code,
		r0 => r0, 
		r1 => r1, 
		r2 => r2, 
		r3 => r3, 
		r4 => r4, 
		r5 => r5, 
		r6 => r6, 
		r7 => r7,
		clk            => clk,
		reset          => reset
	    );
	
	controlpath_risc : controlpath
			port map(
		m_mem_a	       => m_mem_a,
		m_a3_0         => m_a3_0,
		m_a3_1 	       => m_a3_1,
		m_d3_0         => m_d3_0,
		m_d3_1 	       => m_d3_1,
		m_z            => m_z,
		m_op2_0	       => m_op2_0,
		m_op2_1	       => m_op2_1,
		m_a2          => m_a2,
		m_op1_0          => m_op1_0,
		m_op1_1          => m_op1_1,
		wr_mem         => wr_mem,  
		rd_mem         => rd_mem,  
		wr_rf          => wr_rf,   
		en_ir          => en_ir,   
		en_irf      => en_irf, 
		en_A           => en_A,  
		en_c           => en_c,
		m_comp_a       => m_comp_a,
		m_comp_b       => m_comp_b,
		en_z           => en_z,
		op_sel         => op_sel,   
		equ            => equ,    
		C              => C,
		Z              => Z,  
		op_code        => op_code,
		condition_code => condition_code,
		clk            => clk,
		reset          => reset
	    );
		 
		
end behave;
